`include "define.vh"

module alu(
    input reg [5:0] code;
    input reg [31:0] op1;
    input reg [31:0] op2;
    output wire [31:0]  result;
    output wire br;
    );

    always @(*) begin
    
    end

endmodule