module pc (clk)